BZh91AY&SY3r�> F߀Py����װ����P�k����ţZ%=Mf�j��=6��h����a= jz4!5S� hd�    $ԄH'���hdh�� h ��h`LM&L�LM2100	"#B�	��5O$ؓzP  h h�!�ْB��b3��� u�Q���H�4�>�W��L�C�&L����щ�rp�333q�ה���I��wM�Ƃ7��8bw���H�݉}�:����x*�y��x@`�a$`OB�Ⱥ�,+":#]�,E�B��hEa!�_;hj9r�� �G�G?�.��I��S��j1$5n�3~`���J�a�6l0@�e��wN�pX�b&s�!���&�sQJD>��
�1�r*pa*��7�9�)ZMک�V���SK90�;�p㛇u��k�A�݆���3��A�P��rM�9�ML�{��#t��7�ֶ.�%�Dk0a�Nb�q�8(�/�UP`Q���	Fg%ao.@��q�5�59D؂$�ܸ4�fxw,�*gk
(��CC���6x�
��9({�>w{旘�Ѳ��Jd�S��!��[��Q�B�5�o븧�jRӿk��#�1�L���F�@7v��5a��z�:7�s)@�q�U�_�yT�`Ƥ��iڿ��Z��lG�nA1y+yQ��u7/y(�Y�n�"1�{9�m��ߣI��9��yv��K����d��3n�ʣ��h؇G�i��UX3�e�-:@�'�3XH�DNu�"C�NU>�]�[�p*Ar8���D3��CWv$�p�$0��9󔘫�,�%�_�)��@H��s��pR7M��%�`�KA���2"pv�fT��Hm8D�\� 4�-ϪT���S�+��I�<�k ��2�=@�(
� k �#�L��ˌ��x�	��x�:s�Nɗ����#��v�(�0w1@m: z��g ��+�ʔ�2�&t3\s(6.l�~��;�U�	���v)��ک@H����&fwr��­��G&7���R$Anky`EQ:*5HE Z�}8�7Vʩ��4$;%I���l����ܑN$ܱO�